library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL; 

entity RAM is
port(
    clk     : in  std_logic; 
    Adress  : in  std_logic_vector(7 downto 0);
    Data_in : in  std_logic_vector(23 downto 0);
    EnRAM   : in  std_logic; 
    RW      : in  std_logic; 
    Data_out: out std_logic_vector(23 downto 0)
);
end RAM;

architecture Behavioral of RAM is

    type RAM_MEMORY is array (0 to 255) of std_logic_vector(23 downto 0);
    -- R1=Contador T (para delay), R2/R3=Delay, R4=Contador H
signal MEMORY: RAM_MEMORY := (
    -- =================================================================
    -- PROGRAMA 1: 17x+25y-w/4 (Inicia en 0)
    -- T FIJO = 2 (Resultado 122 -> T=2)
    -- =================================================================
    
    -- === CÁLCULO ECUACIÓN (PC 0-7) ===
    0 => "00001011" & "00000000" & "11011000",  -- (PC=0) LW R0, [W] (Offset=216 -> 0+1+216=217)
    1 => "00001011" & "00000001" & "11011000",  -- (PC=1) LW R1, [X] (Offset=216 -> 1+1+216=218)
    2 => "00001011" & "00000010" & "11011000",  -- (PC=2) LW R2, [Y] (Offset=216 -> 2+1+216=219)
    3 => "00011101" & "00000001" & "00010001",  -- (PC=3) MULI R1, 17 
    4 => "00011101" & "00000010" & "00011001",  -- (PC=4) MULI R2, 25 
    5 => "00011110" & "00000000" & "00000100",  -- (PC=5) DIVI R0, 4 
    6 => "00000000" & "00000001" & "00000010",  -- (PC=6) ADD R1, R2 
    7 => "00000001" & "00000001" & "00000000",  -- (PC=7) SUB R1, R0 (R1 = 122)
    
    -- === DISPLAY Y CONTADOR (PC 8-36) ===
    8 => "00100101" & "00000001" & "00000000",  -- (PC=8) DISP R1 (Muestra 122)
    
    -- (INICIO BLOQUE DELAY 10s)
    9 => "00001011" & "00000001" & "11101100",  -- (PC=9) LW R1, [I_VALUE_10S] (Offset=236 -> 9+1+236=246)
    10 => "00001011" & "00000010" & "11101100", -- (PC=10) ETIQUETA_I_10S: LW R2, [J_VALUE] (Offset=236 -> 10+1+236=247)
    11 => "00001011" & "00000011" & "11101100", -- (PC=11) ETIQUETA_J_10S: LW R3, [K_VALUE] (Offset=236 -> 11+1+236=248)
    12 => "00011010" & "00000000" & "00000000", -- (PC=12) ETIQUETA_K_10S: NOP
    13 => "00011100" & "00000011" & "00000001", -- (PC=13) SUBI R3, 1
    14 => "00010010" & "00000000" & "11111101", -- (PC=14) BNZ (a PC=12). Offset = -3
    15 => "00011100" & "00000010" & "00000001", -- (PC=15) SUBI R2, 1
    16 => "00010010" & "00000000" & "11111010", -- (PC=16) BNZ (a PC=11). Offset = -6
    17 => "00011100" & "00000001" & "00000001", -- (PC=17) SUBI R1, 1
    18 => "00010010" & "00000000" & "11110111", -- (PC=18) BNZ (a PC=10). Offset = -9
    -- (FIN BLOQUE DELAY 10s)

    -- (INICIO BLOQUE CONTADOR H=1-30)
    19 => "00001011" & "00000100" & "11100110",  -- (PC=19) LW R4, [H_INIT=1] (Offset=230 -> 19+1+230=250)
    20 => "00100101" & "00000100" & "00000000",  -- (PC=20) ETIQUETA_H_LOOP: DISP R4 (Muestra H)
    -- P1 CARGA T=2 (Addr 249)
    21 => "00001011" & "00000001" & "11100011",  -- (PC=21) LW R1, [T_VAL_2] (Offset=227 -> 21+1+227=249)
    22 => "00001011" & "00000010" & "11100000",  -- (PC=22) ETIQUETA_I_T: LW R2, [J_VALUE] (Offset=224 -> 22+1+224=247)
    23 => "00001011" & "00000011" & "11100000",  -- (PC=23) ETIQUETA_J_T: LW R3, [K_VALUE] (Offset=224 -> 23+1+224=248)
    24 => "00011010" & "00000000" & "00000000",  -- (PC=24) ETIQUETA_K_T: NOP
    25 => "00011100" & "00000011" & "00000001",  -- (PC=25) SUBI R3, 1
    26 => "00010010" & "00000000" & "11111101",  -- (PC=26) BNZ (a PC=24). Offset = -3
    27 => "00011100" & "00000010" & "00000001",  -- (PC=27) SUBI R2, 1
    28 => "00010010" & "00000000" & "11111010",  -- (PC=28) BNZ (a PC=23). Offset = -6
    29 => "00011100" & "00000001" & "00000001",  -- (PC=29) SUBI R1, 1 (Decrementa T)
    30 => "00010010" & "00000000" & "11110111",  -- (PC=30) BNZ (a PC=22). Offset = -9
    31 => "00011011" & "00000100" & "00000001",  -- (PC=31) ADDI R4, 1 (H = H+1)
    32 => "00100011" & "00001111" & "00000001",  -- (PC=32) ASRI R15, 1 (LEDs)
    33 => "00011111" & "00000100" & "00011111",  -- (PC=33) CMPI R4, 31 
    34 => "00010010" & "00000000" & "11110001",  -- (PC=34) BNZ (a PC=20). Offset = -15
    35 => "00100100" & "00000000" & "00000000",  -- (PC=35) HALT
    36 => "00100100" & "00000000" & "00000000",  -- (PC=36) HALT (seguridad)
    -- === FIN PROGRAMA 1 ===

    -- =================================================================
    -- PROGRAMA 2: 10x^2 + 30x - z/2 (Inicia en 37)
    -- T FIJO = 3 (Resultado 90 -> T=3)
    -- =================================================================
    
    -- === CÁLCULO ECUACIÓN (PC 37-45) ===
    37 => "00001011" & "00000000" & "10110100",  -- (PC=37) LW R0, [X] (Offset=180 -> 37+1+180=218)
    38 => "00001011" & "00000001" & "10110011",  -- (PC=38) LW R1, [X] (Offset=179 -> 38+1+179=218)
    39 => "00001011" & "00000010" & "10110100",  -- (PC=39) LW R2, [Z] (Offset=180 -> 39+1+180=220)
    40 => "00000010" & "00000000" & "00000000",  -- (PC=40) MUL R0, R0 (X^2)
    41 => "00011101" & "00000000" & "00001010",  -- (PC=41) MULI R0, 10
    42 => "00011101" & "00000001" & "00011110",  -- (PC=42) MULI R1, 30
    43 => "00000000" & "00000000" & "00000001",  -- (PC=43) ADD R0, R1
    44 => "00011110" & "00000010" & "00000010",  -- (PC=44) DIVI R2, 2
    45 => "00000001" & "00000000" & "00000010",  -- (PC=45) SUB R0, R2 (R0 = 90)

    -- === DISPLAY Y CONTADOR (PC 46-73) ===
    46 => "00100101" & "00000000" & "00000000",  -- (PC=46) DISP R0 (Muestra 90)
    
    -- (INICIO BLOQUE DELAY 10s)
    47 => "00001011" & "00000001" & "11000110",  -- (PC=47) LW R1, [I_VALUE_10S] (Offset=198 -> 47+1+198=246)
    48 => "00001011" & "00000010" & "11000110",  -- (PC=48) ETIQUETA_I_10S: LW R2, [J_VALUE] (Offset=198 -> 48+1+198=247)
    49 => "00001011" & "00000011" & "11000110",  -- (PC=49) ETIQUETA_J_10S: LW R3, [K_VALUE] (Offset=198 -> 49+1+198=248)
    50 => "00011010" & "00000000" & "00000000",  -- (PC=50) ETIQUETA_K_10S: NOP
    51 => "00011100" & "00000011" & "00000001",  -- (PC=51) SUBI R3, 1
    52 => "00010010" & "00000000" & "11111101",  -- (PC=52) BNZ (a PC=50). Offset = -3
    53 => "00011100" & "00000010" & "00000001",  -- (PC=53) SUBI R2, 1
    54 => "00010010" & "00000000" & "11111010",  -- (PC=54) BNZ (a PC=49). Offset = -6
    55 => "00011100" & "00000001" & "00000001",  -- (PC=55) SUBI R1, 1
    56 => "00010010" & "00000000" & "11110111",  -- (PC=56) BNZ (a PC=48). Offset = -9
    -- (FIN BLOQUE DELAY 10s)

    -- (INICIO BLOQUE CONTADOR H=1-30)
    57 => "00001011" & "00000100" & "11000000",  -- (PC=57) LW R4, [H_INIT=1] (Offset=192 -> 57+1+192=250)
    58 => "00100101" & "00000100" & "00000000",  -- (PC=58) ETIQUETA_H_LOOP: DISP R4 (Muestra H)
    -- *** CAMBIO: P2 CARGA T=3 (Addr 252) ***
    59 => "00001011" & "00000001" & "11000000",  -- (PC=59) LW R1, [T_VAL_3] (Offset=192 -> 59+1+192=252)
    60 => "00001011" & "00000010" & "10111010",  -- (PC=60) ETIQUETA_I_T: LW R2, [J_VALUE] (Offset=186 -> 60+1+186=247)
    61 => "00001011" & "00000011" & "10111010",  -- (PC=61) ETIQUETA_J_T: LW R3, [K_VALUE] (Offset=186 -> 61+1+186=248)
    62 => "00011010" & "00000000" & "00000000",  -- (PC=62) ETIQUETA_K_T: NOP
    63 => "00011100" & "00000011" & "00000001",  -- (PC=63) SUBI R3, 1
    64 => "00010010" & "00000000" & "11111101",  -- (PC=64) BNZ (a PC=62). Offset = -3
    65 => "00011100" & "00000010" & "00000001",  -- (PC=65) SUBI R2, 1
    66 => "00010010" & "00000000" & "11111010",  -- (PC=66) BNZ (a PC=61). Offset = -6
    67 => "00011100" & "00000001" & "00000001",  -- (PC=67) SUBI R1, 1 (Decrementa T)
    68 => "00010010" & "00000000" & "11110111",  -- (PC=68) BNZ (a PC=60). Offset = -9
    69 => "00011011" & "00000100" & "00000001",  -- (PC=69) ADDI R4, 1 (H = H+1)
    70 => "00100011" & "00001111" & "00000001",  -- (PC=70) ASRI R15, 1 (LEDs)
    71 => "00011111" & "00000100" & "00011111",  -- (PC=71) CMPI R4, 31 
    72 => "00010010" & "00000000" & "11110001",  -- (PC=72) BNZ (a PC=58). Offset = -15
    73 => "00100100" & "00000000" & "00000000",  -- (PC=73) HALT
    -- === FIN PROGRAMA 2 ===

    -- =================================================================
    -- PROGRAMA 3: -X^3 – 7Z+ W / (10) (Inicia en 74)
    -- T FIJO = 5 (Resultado -143 -> T=5)
    -- =================================================================
    
    -- === CÁLCULO ECUACIÓN (PC 74-82) ===
    74 => "00001011" & "00000000" & "10001110",  -- (PC=74) LW R0, [W] (Offset=142 -> 74+1+142=217)
    75 => "00001011" & "00000001" & "10001110",  -- (PC=75) LW R1, [X] (Offset=142 -> 75+1+142=218)
    76 => "00001011" & "00000010" & "10001111",  -- (PC=76) LW R2, [Z] (Offset=143 -> 76+1+143=220)
    77 => "00001011" & "00000011" & "10001100",  -- (PC=77) LW R3, [X] (Offset=140 -> 77+1+140=218)
    78 => "00000010" & "00000001" & "00000001",  -- (PC=78) MUL R1, R1 (X^2)
    79 => "00000010" & "00000001" & "00000011",  -- (PC=79) MUL R1, R3 (X^3)
    80 => "00011101" & "00000010" & "00000111",  -- (PC=80) MULI R2, 7 (7Z)
    81 => "00011110" & "00000000" & "00001010",  -- (PC=81) DIVI R0, 10 (W/10)
    82 => "00000001" & "00000000" & "00000010",  -- (PC=82) SUB R0, R2
    83 => "00000001" & "00000000" & "00000001",  -- (PC=83) SUB R0, R1 (R0 = -143)
    
    -- === DISPLAY Y CONTADOR (PC 84-111) ===
    84 => "00100101" & "00000000" & "00000000",  -- (PC=84) DISP R0 (Muestra -143)
    
    -- (INICIO BLOQUE DELAY 10s)
    85 => "00001011" & "00000001" & "10100000",  -- (PC=85) LW R1, [I_VALUE_10S] (Offset=160 -> 85+1+160=246)
    86 => "00001011" & "00000010" & "10100000",  -- (PC=86) ETIQUETA_I_10S: LW R2, [J_VALUE] (Offset=160 -> 86+1+160=247)
    87 => "00001011" & "00000011" & "10100000",  -- (PC=87) ETIQUETA_J_10S: LW R3, [K_VALUE] (Offset=160 -> 87+1+160=248)
    88 => "00011010" & "00000000" & "00000000",  -- (PC=88) ETIQUETA_K_10S: NOP
    89 => "00011100" & "00000011" & "00000001",  -- (PC=89) SUBI R3, 1
    90 => "00010010" & "00000000" & "11111101",  -- (PC=90) BNZ (a PC=88). Offset = -3
    91 => "00011100" & "00000010" & "00000001",  -- (PC=91) SUBI R2, 1
    92 => "00010010" & "00000000" & "11111010",  -- (PC=92) BNZ (a PC=87). Offset = -6
    93 => "00011100" & "00000001" & "00000001",  -- (PC=93) SUBI R1, 1
    94 => "00010010" & "00000000" & "11110111",  -- (PC=94) BNZ (a PC=86). Offset = -9
    -- (FIN BLOQUE DELAY 10s)

    -- (INICIO BLOQUE CONTADOR H=1-30)
    95 => "00001011" & "00000100" & "10011010",  -- (PC=95) LW R4, [H_INIT=1] (Offset=154 -> 95+1+154=250)
    96 => "00100101" & "00000100" & "00000000",  -- (PC=96) ETIQUETA_H_LOOP: DISP R4 (Muestra H)
    -- *** CAMBIO: P3 CARGA T=5 (Addr 254) ***
    97 => "00001011" & "00000001" & "10011100",  -- (PC=97) LW R1, [T_VAL_5] (Offset=156 -> 97+1+156=254)
    98 => "00001011" & "00000010" & "10010100",  -- (PC=98) ETIQUETA_I_T: LW R2, [J_VALUE] (Offset=148 -> 98+1+148=247)
    99 => "00001011" & "00000011" & "10010100",  -- (PC=99) ETIQUETA_J_T: LW R3, [K_VALUE] (Offset=148 -> 99+1+148=248)
    100 => "00011010" & "00000000" & "00000000", -- (PC=100) ETIQUETA_K_T: NOP
    101 => "00011100" & "00000011" & "00000001", -- (PC=101) SUBI R3, 1
    102 => "00010010" & "00000000" & "11111101", -- (PC=102) BNZ (a PC=100). Offset = -3
    103 => "00011100" & "00000010" & "00000001", -- (PC=103) SUBI R2, 1
    104 => "00010010" & "00000000" & "11111010", -- (PC=104) BNZ (a PC=99). Offset = -6
    105 => "00011100" & "00000001" & "00000001", -- (PC=105) SUBI R1, 1 (Decrementa T)
    106 => "00010010" & "00000000" & "11110111", -- (PC=106) BNZ (a PC=98). Offset = -9
    107 => "00011011" & "00000100" & "00000001", -- (PC=107) ADDI R4, 1 (H = H+1)
    108 => "00100011" & "00001111" & "00000001", -- (PC=108) ASRI R15, 1 (LEDs)
    109 => "00011111" & "00000100" & "00011111", -- (PC=109) CMPI R4, 31 
    110 => "00010010" & "00000000" & "11110001", -- (PC=110) BNZ (a PC=96). Offset = -15
    111 => "00100100" & "00000000" & "00000000", -- (PC=111) HALT
    -- === FIN PROGRAMA 3 ===

    -- =================================================================
    -- PROGRAMA 4: HALT (Inicia en 112)
    -- =================================================================
    112 => "00100100" & "00000000" & "00000000",  -- (PC=112) HALT
    -- === FIN PROGRAMA 4 ===


    -- =================================================================
    -- SECCIÓN DE DATOS
    -- =================================================================
    -- *** NUEVOS VALORES W,X,Y,Z ***
    217 => "00000000" & "00000000" & "00110010",  -- W = 50 decimal
    218 => "00000000" & "00000000" & "00000010",  -- X = 2 decimal
    219 => "00000000" & "00000000" & "00000100",  -- Y = 4 decimal
    220 => "00000000" & "00000000" & "00010100",  -- Z = 20 decimal
    
    -- Constantes de Delays (Reutilizadas)
    246 => "00000000" & "00000000" & "00001010",  -- I_VALUE_10S = 10
    247 => "00000000" & "00000000" & "00100101",  -- J_VALUE = 37
    248 => "00000000" & "11111111" & "11111111",  -- K_VALUE = 65535

    -- Constantes para T y H (Contador 1-30)
    249 => "00000000" & "00000000" & "00000010",  -- T_VAL_2 (para P1)
    250 => "00000000" & "00000000" & "00000001",  -- H_INIT = 1
    
    -- *** DATOS T AÑADIDOS ***
    251 => "00000000" & "00000000" & "00000001",  -- T_VAL_1 = 1
    252 => "00000000" & "00000000" & "00000011",  -- T_VAL_3 (para P2)
    253 => "00000000" & "00000000" & "00000100",  -- T_VAL_4 = 4
    254 => "00000000" & "00000000" & "00000101",  -- T_VAL_5 (para P3)
    

    others => (others => '0')
);
    
    signal addr_int : integer range 0 to 255; 
--    
begin
 
    addr_int <= to_integer(unsigned(Adress));
 
    -- Escritura Síncrona
    process(clk)
    begin
        if rising_edge(clk) then
            if EnRAM = '1' and RW = '0' then 
                MEMORY(addr_int) <= Data_in;
            end if;
        end if;
    end process;

    -- Lectura Asíncrona
    Data_out <= MEMORY(addr_int);

end Behavioral;